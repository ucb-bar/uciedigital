`timescale 1ps/1ps

// Positive edge triggered D flip-flop
module pos_dff #(
    parameter real T_CLKQ = 5.0   // Clock-to-q delay in ps
)(
    input logic clk,
    input logic d,
    input logic rstb,
    output logic q
);

    specify
        specparam T_SETUP = 5.0;  // Setup time in ps
        specparam T_HOLD = 2.0;  // Hold time in ps
        $setup(d, posedge clk, T_SETUP);
        $hold(posedge clk, d, T_HOLD);
    endspecify

    // TODO: design reset distribution/async reset?
    always_ff @(posedge clk, negedge rstb) begin
        if (!rstb)
            q <= 1'b0;
        else
            q <= #(T_CLKQ) d;
    end
endmodule


module tb_dff;

    // Signals
    logic clk;
    logic d;
    logic q;

    // Ips DUT
    pos_dff #(
        .T_CLKQ(5.0)
    ) dut (
        .clk(clk),
        .d(d),
        .q(q)
    );

    // Clock generation (10ps period)
    initial clk = 0;
    always #5 clk = ~clk;

    // Test stimulus
    initial begin
        d = 0;

        repeat (2) @(posedge clk);

        // --- Setup violation: change 'd' too close to clock ---
        $display("Testing setup violation at %0t", $time);
        #7 // 3ps before clk edge, setup required is 5ps
        d = 1;
        @(posedge clk);

        repeat (2) @(posedge clk);

        // --- Hold violation: change 'd' too soon after clock ---
        $display("Testing hold violation at %0t", $time);
        @(posedge clk);
        #1;  // 1ps after clk edge, hold required is 2ps
        d = 0;

        repeat (2) @(posedge clk);

        // Normal operation (no violation)
        $display("Normal operation at %0t", $time);
        @(posedge clk);
        #3 // 3ps after clk edge and 7ps before next clk edge, satisfies setup/hold
        d = 1;
        @(posedge clk);
        #6 // Wait for data-to-q delay.
        if (q != 1'b1) $error("Incorrect q value (expected %b, got %b)", d, q);
        @(posedge clk);
        #3
        d = 0;
        @(posedge clk);
        #6
        if (q != 1'b0) $error("Incorrect q value (expected %b, got %b)", d, q);

        repeat (2) @(posedge clk);

        $finish;
    end

endmodule

// Positive transparent latch
module pos_latch #(
    parameter real T_CLKQ_DQ = 5.0     // Clock-to-q and data-to-q delay in ps.
)(
    input logic clk,
    input logic d,
    output logic q
);

    specify
        specparam T_SETUP = 5.0;  // Setup time in ps
        specparam T_HOLD  = 2.0;  // Hold time in ps
        $setup(d, negedge clk, T_SETUP);
        $hold(negedge clk, d, T_HOLD);
    endspecify

    always_latch begin
        if (clk) begin
            q <= #(T_CLKQ_DQ) d;
        end
    end
endmodule

// Negative transparent latch
module neg_latch #(
    parameter real T_CLKQ_DQ = 5.0     // Clock-to-q and data-to-q delay in ps.
)(
    input logic clkb,
    input logic d,
    output logic q
);

    specify
        specparam T_SETUP = 5.0;  // Setup time in ps
        specparam T_HOLD  = 2.0;  // Hold time in ps
        $setup(d, posedge clkb, T_SETUP);
        $hold(posedge clkb, d, T_HOLD);
    endspecify

    always_latch begin
        if (!clkb) begin
            q <= #(T_CLKQ_DQ) d;
        end
    end
endmodule


module tb_latch;

    logic clk;
    logic clkb;
    logic d;
    logic qp;
    logic qn;

    pos_latch #(
        .T_CLKQ_DQ(5.0)
    ) pdut (
        .clk(clk),
        .d(d),
        .q(qp)
    );

    neg_latch #(
        .T_CLKQ_DQ(5.0)
    ) ndut (
        .clkb(clkb),
        .d(d),
        .q(qn)
    );

    // Clock generation (10ps period)
    initial clk = 0;
    always #5 clk = ~clk;
    assign clkb = ~clk;

    // Test stimulus
    initial begin
        d = 0;

        // Negedge is the sampling edge for positive transparent latches.
        repeat (2) @(negedge clk);

        // --- Setup violation: change 'd' too close to clock ---
        $display("Testing setup violation at %0t", $time);
        #8 // 2ps before clk edge, setup required is 5ps
        d = 1;

        repeat (2) @(negedge clk);

        // --- Hold violation: change 'd' too soon after clock ---
        $display("Testing hold violation at %0t", $time);
        @(negedge clk);
        #1;  // 1ps after clk edge, hold required is 2ps
        d = 0;

        repeat (2) @(negedge clk);

        // Normal operation (no violation)
        $display("Normal operation at %0t", $time);
        @(negedge clk);
        #3 // 3ps after clk edge and 7ps before next clk edge, satisfies setup/hold
        d = 1;
        @(negedge clk);
        #6 // Output should be up after T_CLKQ_DQ delay.
        if (qp != 1'b1) $error("Incorrect q value for pos_latch (expected %b, got %b)", d, qp);
        if (qn != 1'b1) $error("Incorrect q value for neg_latch (expected %b, got %b)", d, qn);
        @(negedge clk);
        #3
        d = 0;
        @(negedge clk);
        #6
        if (qp != 1'b0) $error("Incorrect q value for pos_latch (expected %b, got %b)", d, qp);
        if (qn != 1'b0) $error("Incorrect q value for neg_latch (expected %b, got %b)", d, qn);

        repeat (2) @(negedge clk);

        $finish;
    end

endmodule

module mux #(
    parameter real DELAY = 5.0 // Delay in ps.
)(
    input logic sel_a,
    input logic a,
    input logic b,
    output logic o
);
    assign #(DELAY) o = sel_a ? a : b;
endmodule
